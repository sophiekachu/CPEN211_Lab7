module vDFFE(clk, load, in, out) ;
  parameter n = 16;  // width
  input clk, load ;
  input  [n-1:0] in ;
  output [n-1:0] out ;
  reg    [n-1:0] out ;
  wire   [n-1:0] next_out;

  assign next_out = load ? in : out;

  always @(posedge clk)
    out = next_out;
endmodule 
